interface uart_if;

  logic RXD;
  logic TXD;

endinterface: uart_if
